module tb_fixedpoint_formatter ();
    
parameter WIDTH_INPUT       = 32;
parameter WIDTH_OUTPUT      = 16;
parameter WIDTH_INTEGER     = 6 ;
parameter WIDTH_FRACTION    = 9 ;

logic   [WIDTH_INPUT - 1 : 0]   data_i;
logic   [WIDTH_OUTPUT - 1 : 0]  data_o; 

fixedpoint_formatter #(
    .WIDTH_INPUT(WIDTH_INPUT),
    .WIDTH_OUTPUT(WIDTH_OUTPUT),
    .WIDTH_INTEGER(WIDTH_INTEGER),
    .WIDTH_FRACTION(WIDTH_FRACTION)
) fixedpoint_formatter_inst (
    .data_i(data_i),
    .data_o(data_o)
);

initial begin
    $dumpfile("./out/tb_fixedpoint_formatter.vcd");
    $dumpvars(0, tb_fixedpoint_formatter);
end

initial begin
    // pos
    data_i = 32'b00000000_000000_000000000_000000000;
    #10;
    data_i = 32'b00000000_000000_000000000_100000000;
    #10;
    data_i = 32'b00000000_000000_000000001_100000000;
    #10;
    data_i = 32'b00000000_000000_111111111_100000000;
    #10;
    data_i = 32'b00000000_000000_000000000_010000000;
    #10;
    data_i = 32'b00000000_000000_000000001_010000000;
    #10;
    data_i = 32'b00000000_000000_111111111_010000000;
    #10;
    // pos sat
    data_i = 32'b00000001_000000_000000000_000000000;
    #10;
    data_i = 32'b00000001_000000_000000000_100000000;
    #10;
    data_i = 32'b00000001_000000_000000001_100000000;
    #10;
    data_i = 32'b00000001_000000_111111111_100000000;
    #10;
    data_i = 32'b00000001_000000_000000000_010000000;
    #10;
    data_i = 32'b00000001_000000_000000001_010000000;
    #10;
    data_i = 32'b00000001_000000_111111111_010000000;
    #10;

    // neg
    data_i = 32'b11111111_000000_000000000_000000000;
    #10;
    data_i = 32'b11111111_000000_000000000_100000000;
    #10;
    data_i = 32'b11111111_000000_000000000_110000000;
    #10;
    data_i = 32'b11111111_100000_000000000_000000000;
    #10;
    data_i = 32'b11111111_100000_000000000_100000000;
    #10;
    data_i = 32'b11111111_100000_000000000_101000000;
    #10;
    data_i = 32'b11111111_100000_000000001_100000000;
    #10;
    data_i = 32'b11111111_100000_000000001_101000000;
    #10;
    data_i = 32'b11111111_111111_111111111_100000000;
    #10;
    data_i = 32'b11111111_111111_111111111_100010000;
    #10;
    data_i = 32'b11111111_111111_111111111_010000000;
    #10;
    data_i = 32'b11111111_111111_111111111_010010000;
    #10;

    // neg sat
    data_i = 32'b11011111_000000_000000000_000000000;
    #10;
    data_i = 32'b11011111_000000_000000000_100000000;
    #10;
    data_i = 32'b11011111_000000_000000000_110000000;
    #10;
    data_i = 32'b11011111_100000_000000000_000000000;
    #10;
    data_i = 32'b11011111_100000_000000000_100000000;
    #10;
    data_i = 32'b11011111_100000_000000000_101000000;
    #10;
    data_i = 32'b11011111_100000_000000001_100000000;
    #10;
    data_i = 32'b11011111_100000_000000001_101000000;
    #10;
    data_i = 32'b11011111_111111_111111111_100000000;
    #10;
    data_i = 32'b11011111_111111_111111111_100010000;
    #10;
    data_i = 32'b11011111_111111_111111111_010000000;
    #10;
    data_i = 32'b11011111_111111_111111111_010010000;
    #10;

    data_i = 32'b00000000_000000_000000000_000000000;
    #10;
end

endmodule