///////////////////////////////////////////////////////////
// Author: Jackbang
///////////////////////////////////////////////////////////

